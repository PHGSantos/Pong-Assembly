	component nios is
		port (
			btn_external_connection_export : in  std_logic                    := 'X'; -- export
			clk_clk                        : in  std_logic                    := 'X'; -- clk
			led_external_connection_export : out std_logic_vector(7 downto 0);        -- export
			reset_reset_n                  : in  std_logic                    := 'X'  -- reset_n
		);
	end component nios;

	u0 : component nios
		port map (
			btn_external_connection_export => CONNECTED_TO_btn_external_connection_export, -- btn_external_connection.export
			clk_clk                        => CONNECTED_TO_clk_clk,                        --                     clk.clk
			led_external_connection_export => CONNECTED_TO_led_external_connection_export, -- led_external_connection.export
			reset_reset_n                  => CONNECTED_TO_reset_reset_n                   --                   reset.reset_n
		);

